module endpoint_ctrl (
	input NRST,
	input CLK,
	input [23:0] TOKEN_IN,
	input TOKEN_IN_STRB,
	input [7:0] DATA_IN,
	input DATA_IN_STRB,
	input DATA_IN_END,
	input DATA_IN_FAIL
);

endmodule
